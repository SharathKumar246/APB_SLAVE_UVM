package apb_pkg;
import uvm_pkg::*;
`include "uvm_macros.svh"
  `include "apb_sequence_item.sv"
  `include "apb_sequence.sv"
  `include "apb_sequencer.sv"
  `include "apb_driver.sv"
  `include "apb_active_monitor.sv"
  `include "apb_passive_monitor.sv"
  `include "apb_active_agent.sv"
  `include "apb_passive_agent.sv"
  `include "apb_scoreboard.sv"
  `include "apb_subscriber.sv"
  `include "apb_environment.sv"
  `include "apb_test.sv"

endpackage